module control(input Run, ClearA_LoadB, Reset, output Clr_Ld, Shift, Add, Sub);
