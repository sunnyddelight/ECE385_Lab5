module computation_module(input [8:0] A, B,
							input Add, Sub, Clr_Ld,
							output[8:0] S);

						assign S=A;
							
endmodule
